-- include libraries
-- standard stuff
library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

PACKAGE PromPkg IS
END PromPkg;

PACKAGE BODY PromPkg IS
END PromPkg;

library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Prom is
  GENERIC(
    addr_width : integer := 16384; -- store 128 elements (512 bytes)
    addr_bits  : integer := 14; -- required bits to store 128 elements
    data_width : integer := 32 -- each element has 32-bits
    );
  PORT(
    addr : IN std_logic_vector(addr_bits-1 downto 0);
    data : OUT std_logic_vector(data_width-1 downto 0)
    );
end Prom;

architecture arch of Prom is

  type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);
  
  signal Prom_ROM : rom_type := (
-- copy/paste the ROM content here --
"11110001000010000100100001000000", -- 1
"00000000000000000000000100011100", -- 2
"00010010000011010101001001000100", -- 3
"01001111010011000010110001010011", -- 4
"01000010011101010111001101000110", -- 5
"01010000010001110100000100000010", -- 6
"00000001000000010000001000010000", -- 7
"00000000000000010000000000000000", -- 8
"00011110000000010000001100010000", -- 9
"00000000000000000000000100000000", -- 10
"00000001000101100001000000000000", -- 11
"00000000000000000111111100000001", -- 12
"00010001000100100001000101110011", -- 13
"01101100011000010111011001100101", -- 14
"00101101011000100111010101110010", -- 15
"01110011011101000010110101110011", -- 16
"01101001011110100110010101110011", -- 17
"00000001000100000001000000000000", -- 18
"00000000000000000111111100000001", -- 19
"00010001000100100000101101100010", -- 20
"01110101011100100111001101110100", -- 21
"00101101011100110110100101111010", -- 22
"01100101011100110000000100010000", -- 23
"10100100110000001011011000001000", -- 24
"01101100011001010110010000101101", -- 25
"01110110011010010111001001110100", -- 26
"00001000000000001011100000000001", -- 27
"00000010101101100000111101101101", -- 28
"01111001001011010111001101100010", -- 29
"01110101011100110010110101100001", -- 30
"01100100011001000111001001100101", -- 31
"01110011011100110000100000000001", -- 32
"10111010000000010000001110110110", -- 33
"00001101011011010111100100101101", -- 34
"01110011011000100111010101110011", -- 35
"00101101011100110111000001100001", -- 36
"01100011011001010000100000000010", -- 37
"10111010101101100000011001101101", -- 38
"01100001011100000010110101101001", -- 39
"01101110000010000000001110110111", -- 40
"00010010000001100110110101100001", -- 41
"01110000001011010110100101101110", -- 42
"00000010000010011100001010110110", -- 43
"00000111011011010110000101110000", -- 44
"00101101011011110111010101110100", -- 45
"00001000000001001011011100010010", -- 46
"00000111011011010110000101110000", -- 47
"00101101011011110111010101110100", -- 48
"00000010000010011100001010110110", -- 49
"00001010011011010110000101110000", -- 50
"00101101011010010110111000101101", -- 51
"01101100011001010110010000001000", -- 52
"00000101101101110000100000000001", -- 53
"00010000000000000000000100000000", -- 54
"00000000000111100000100000000010", -- 55
"00010000000000000000000000000000", -- 56
"00000100000010000000001111000011", -- 57
"00001000000000001100001010110110", -- 58
"00001011011011010110000101110000", -- 59
"00101101011011110111010101110100", -- 60
"00101101011011000110010101100100", -- 61
"00001000000001101011011100001000", -- 62
"00000000000100000000000000000000", -- 63
"00000000000001000000100000000100", -- 64
"11000010110010100000011001100010", -- 65
"01101100011010010110111001101011", -- 66
"00100001000010000000011110110111", -- 67
"00001000000001010000100000000000", -- 68
"01110011000010000000011011000010", -- 69
"00010000101000000101000000001010", -- 70
"00000101000010000000011100000000", -- 71
-- ROM then filled with zero
    others => (others => '0'));
begin
  data <= Prom_ROM(conv_integer(unsigned(addr)));
end arch; 
