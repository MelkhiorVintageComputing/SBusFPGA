-- include libraries
-- standard stuff
library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

PACKAGE PromPkg IS
END PromPkg;

PACKAGE BODY PromPkg IS
END PromPkg;

library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Prom is
  GENERIC(
    addr_width : integer := 16384; -- store 128 elements (512 bytes)
    addr_bits  : integer := 14; -- required bits to store 128 elements
    data_width : integer := 32 -- each element has 32-bits
    );
  PORT(
    addr : IN std_logic_vector(addr_bits-1 downto 0);
    data : OUT std_logic_vector(data_width-1 downto 0)
    );
end Prom;

architecture arch of Prom is

  type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);

  signal Prom_ROM : rom_type := (
-- copy/paste the ROM content here --
"11110001000010001010010100101001", -- 1
"00000000000000000000001001111010", -- 2
"00010010000100010101001001000100", -- 3
"01001111010011000010110001100011", -- 4
"01110010011110010111000001110100", -- 5
"01101111011001010110111001100111", -- 6
"01101001011011100110010100000010", -- 7
"00000001000000010000001000010000", -- 8
"00000000000000010000000000000000", -- 9
"00011110000000010000001100010000", -- 10
"00000000000000000000000100000000", -- 11
"00000001000101100001000000000000", -- 12
"00000000000000000111111100000001", -- 13
"00010001000100100001000101110011", -- 14
"01101100011000010111011001100101", -- 15
"00101101011000100111010101110010", -- 16
"01110011011101000010110101110011", -- 17
"01101001011110100110010101110011", -- 18
"00000001000100000001000000000000", -- 19
"00000000000000000111111100000001", -- 20
"00010001000100100000101101100010", -- 21
"01110101011100100111001101110100", -- 22
"00101101011100110110100101111010", -- 23
"01100101011100110000000100010000", -- 24
"10100100110000001011011000001000", -- 25
"01101100011001010110010000101101", -- 26
"01110110011010010111001001110100", -- 27
"00001000000000001011100000000001", -- 28
"00000010101101100000111101101101", -- 29
"01111001001011010111001101100010", -- 30
"01110101011100110010110101100001", -- 31
"01100100011001000111001001100101", -- 32
"01110011011100110000100000000001", -- 33
"10111010000000010000001110110110", -- 34
"00001101011011010111100100101101", -- 35
"01110011011000100111010101110011", -- 36
"00101101011100110111000001100001", -- 37
"01100011011001010000100000000010", -- 38
"10111010101101100000011001101101", -- 39
"01100001011100000010110101101001", -- 40
"01101110000010000000001110110111", -- 41
"00010010000001100110110101100001", -- 42
"01110000001011010110100101101110", -- 43
"00000010000010011100001010110110", -- 44
"00000111011011010110000101110000", -- 45
"00101101011011110111010101110100", -- 46
"00001000000001001011011100010010", -- 47
"00000111011011010110000101110000", -- 48
"00101101011011110111010101110100", -- 49
"00000010000010011100001010110110", -- 50
"00001010011011010110000101110000", -- 51
"00101101011010010110111000101101", -- 52
"01101100011001010110010000001000", -- 53
"00000101101101110000100000000001", -- 54
"00010000000000000000000100000000", -- 55
"00000000000111100000100000000010", -- 56
"00010000000000000000000000000000", -- 57
"00000100000010000000001111000011", -- 58
"00001000000000001100001010110110", -- 59
"00001011011011010110000101110000", -- 60
"00101101011011110111010101110100", -- 61
"00101101011011000110010101100100", -- 62
"00001000000001101011011100001000", -- 63
"00000000000100000000000000000000", -- 64
"00000000000001000000100000000100", -- 65
"11000010101101100000011001100010", -- 66
"01101100011010010110111001101011", -- 67
"00100001000010000000011110110111", -- 68
"00001000000001010000100000000000", -- 69
"01110011000010000000011011000010", -- 70
"00010000101000000101000000001010", -- 71
"00000101000010000000011100000001", -- 72
"00100111000000010001111100010010", -- 73
"00001001010100100100010001001111", -- 74
"01001100001011000111010001110010", -- 75
"01101110011001110000001000000001", -- 76
"00000001000000100001000000000000", -- 77
"00000010000000000000000000011110", -- 78
"00000001000000110001000000000000", -- 79
"00000000000000010000000000000001", -- 80
"00010110000100000000000000000000", -- 81
"00000000000001000000000100010001", -- 82
"00010010000100010111001101101100", -- 83
"01100001011101100110010100101101", -- 84
"01100010011101010111001001110011", -- 85
"01110100001011010111001101101001", -- 86
"01111010011001010111001100000001", -- 87
"00010000000100000000000000000000", -- 88
"00000000000001000000000100010001", -- 89
"00010010000010110110001001110101", -- 90
"01110010011100110111010000101101", -- 91
"01110011011010010111101001100101", -- 92
"01110011000000010001000000000001", -- 93
"00000010101101100000111101101101", -- 94
"01111001001011010111001101100010", -- 95
"01110101011100110010110101100001", -- 96
"01100100011001000111001001100101", -- 97
"01110011011100110000100000001000", -- 98
"10111010000000010000001110110110", -- 99
"00001101011011010111100100101101", -- 100
"01110011011000100111010101110011", -- 101
"00101101011100110111000001100001", -- 102
"01100011011001010000100000001001", -- 103
"10111010101101100000011001101101", -- 104
"01100001011100000010110101101001", -- 105
"01101110000010000000101010110111", -- 106
"00010010000001100110110101100001", -- 107
"01110000001011010110100101101110", -- 108
"00000010000010011100001010110110", -- 109
"00000111011011010110000101110000", -- 110
"00101101011011110111010101110100", -- 111
"00001000000010111011011100010010", -- 112
"00000111011011010110000101110000", -- 113
"00101101011011110111010101110100", -- 114
"00000010000010011100001000000001", -- 115
"00100111000000010001111100010010", -- 116
"00001011010100100100010001001111", -- 117
"01001100001011000111001101100100", -- 118
"01100011011000010111001001100100", -- 119
"00000010000000010000000100000010", -- 120
"00010000000000000000001100000000", -- 121
"00000000000111100000000100000011", -- 122
"00010000000000000000000000000001", -- 123
"00000000000000010001011000010000", -- 124
"00000000000000000000000000000100", -- 125
"00000001000100010001001000010001", -- 126
"01110011011011000110000101110110", -- 127
"01100101001011010110001001110101", -- 128
"01110010011100110111010000101101", -- 129
"01110011011010010111101001100101", -- 130
"01110011000000010001000000010000", -- 131
"00000000000000000000000000000100", -- 132
"00000001000100010001001000001011", -- 133
"01100010011101010111001001110011", -- 134
"01110100001011010111001101101001", -- 135
"01111010011001010111001100000001", -- 136
"00010000000000010000001010110110", -- 137
"00001111011011010111100100101101", -- 138
"01110011011000100111010101110011", -- 139
"00101101011000010110010001100100", -- 140
"01110010011001010111001101110011", -- 141
"00001000000011001011101000000001", -- 142
"00000011101101100000110101101101", -- 143
"01111001001011010111001101100010", -- 144
"01110101011100110010110101110011", -- 145
"01110000011000010110001101100101", -- 146
"00001000000011011011101010110110", -- 147
"00000110011011010110000101110000", -- 148
"00101101011010010110111000001000", -- 149
"00001110101101110001001000000110", -- 150
"01101101011000010111000000101101", -- 151
"01101001011011100000001000001001", -- 152
"11000010101101100000011101101101", -- 153
"01100001011100000010110101101111", -- 154
"01110101011101000000100000001111", -- 155
"10110111000100100000011101101101", -- 156
"01100001011100000010110101101111", -- 157
"01110101011101000000001000001001", -- 158
"11000010000000000000000000000000", -- 159
-- ROM then filled with zero
    others => (others => '0'));
begin
  data <= Prom_ROM(conv_integer(unsigned(addr)));
end arch; 
