-- include libraries
-- standard stuff
library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

PACKAGE PromPkg IS
END PromPkg;

PACKAGE BODY PromPkg IS
END PromPkg;

library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Prom is
  GENERIC(
    addr_width : integer := 128; -- store 128 elements (512 bytes)
    addr_bits  : integer := 7; -- required bits to store 128 elements
    data_width : integer := 32 -- each element has 32-bits
    );
  PORT(
    addr : IN std_logic_vector(addr_bits-1 downto 0);
    data : OUT std_logic_vector(data_width-1 downto 0)
    );
end Prom;

architecture arch of Prom is

  type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);
  
  signal Prom_ROM : rom_type := (
-- copy/paste the ROM content here --
"11111101000010000000010001111001", -- 1
"00000000000000000000000000101011", -- 2
"00010010000011010101001001000100", -- 3
"01001111010011000010110001010011", -- 4
"01000010011101010111001101000110", -- 5
"01010000010001110100000100000010", -- 6
"00000001000000010000001000010000", -- 7
"00000000000000000000001000000000", -- 8
"00011110000000010000001100010000", -- 9
"00000000000000000000000100000000", -- 10
"00000001000101100000000000000000", -- 11

--    "11111101000010000001001000110001", -- 1
--    "00000000000000000000000001100001", -- 2
--    "10000111000100100000110101010010", -- 3
--    "01000100010011110100110000101100", -- 4
--    "01010011010000100111010101110011", -- 5
--    "01000110010100000100011101000001", -- 6
--    "00000001000101000001001000000100", -- 7
--    "01101110011000010110110101100101", -- 8
--    "00000001000100000000000100000010", -- 9
--    "00010000000000000000000000000010", -- 10
--    "00000000000111100000000100000011", -- 11
--    "00010000000000000000000000000000", -- 12
--    "00000100000100100000001101110010", -- 13
--    "01100101011001110000000100010000", -- 14
--    "00010000000000000000000000000000", -- 15
--    "00010101000100100001000101110011", -- 16
--    "01101100011000010111011001100101", -- 17
--    "00101101011000100111010101110010", -- 18
--    "01110011011101000010110101110011", -- 19
--    "01101001011110100110010101110011", -- 20
--    "00000001000100001011010100001000", -- 21
--    "00000000101101110000000100000010", -- 22
--    "00010000000000000000000000000010", -- 23
--    "00000000000111100111001011000010", -- 24
-- ROM then filled with zero
    others => (others => '0'));
begin
  data <= Prom_ROM(conv_integer(unsigned(addr)));
end arch; 
