-- include libraries
-- standard stuff
library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

PACKAGE PromPkg IS
END PromPkg;

PACKAGE BODY PromPkg IS
END PromPkg;

library IEEE;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Prom is
  GENERIC(
    addr_width : integer := 128; -- store 128 elements (512 bytes)
    addr_bits  : integer := 7; -- required bits to store 128 elements
    data_width : integer := 32 -- each element has 32-bits
    );
  PORT(
    addr : IN std_logic_vector(addr_bits-1 downto 0);
    data : OUT std_logic_vector(data_width-1 downto 0)
    );
end Prom;

architecture arch of Prom is

  type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);
  
  signal Prom_ROM : rom_type := (
-- copy/paste the ROM content here --
"11110001000010000100001101110100", -- 1
"00000000000000000000000100000110", -- 2
"00010010000011010101001001000100", -- 3
"01001111010011000010110001010011", -- 4
"01000010011101010111001101000110", -- 5
"01010000010001110100000100000010", -- 6
"00000001000000010000001000010000", -- 7
"00000000000000000000001000000000", -- 8
"00011110000000010000001100010000", -- 9
"00000000000000000000000100000000", -- 10
"00000001000101100001000000000000", -- 11
"00000000000000000111111100000001", -- 12
"00010001000100100001000101110011", -- 13
"01101100011000010111011001100101", -- 14
"00101101011000100111010101110010", -- 15
"01110011011101000010110101110011", -- 16
"01101001011110100110010101110011", -- 17
"00000001000100001010010011000000", -- 18
"11001010000010000110110001100101", -- 19
"01100100001011010111011001101001", -- 20
"01110010011101000000100000000000", -- 21
"10111000000000010000001011001010", -- 22
"00001111011011010111100100101101", -- 23
"01110011011000100111010101110011", -- 24
"00101101011000010110010001100100", -- 25
"01110010011001010111001101110011", -- 26
"00001000000000011011101000000001", -- 27
"00000011110010100000110101101101", -- 28
"01111001001011010111001101100010", -- 29
"01110101011100110010110101110011", -- 30
"01110000011000010110001101100101", -- 31
"00001000000000101011101011001010", -- 32
"00000110011011010110000101110000", -- 33
"00101101011010010110111000001000", -- 34
"00000011101101110001001000000110", -- 35
"01101101011000010111000000101101", -- 36
"01101001011011100000001000001001", -- 37
"11000010110010100000011101101101", -- 38
"01100001011100000010110101101111", -- 39
"01110101011101000000100000000100", -- 40
"10110111000100100000011101101101", -- 41
"01100001011100000010110101101111", -- 42
"01110101011101000000001000001001", -- 43
"11000010110010100000101001101101", -- 44
"01100001011100000010110101101001", -- 45
"01101110001011010110110001100101", -- 46
"01100100000010000000010110110111", -- 47
"00001000000000010001000000000000", -- 48
"00000000000000100000000000011110", -- 49
"00001000000000100001000000000000", -- 50
"00000000000000000000010000001000", -- 51
"00000011110000110000100000000000", -- 52
"11000010110010100000101101101101", -- 53
"01100001011100000010110101101111", -- 54
"01110101011101000010110101101100", -- 55
"01100101011001000000100000000110", -- 56
"10110111000010000000000000010000", -- 57
"00000000000000000000000000000100", -- 58
"00001000000001001100001011001010", -- 59
"00000110011000100110110001101001", -- 60
"01101110011010110010000100001000", -- 61
"00000111101101110000100000000101", -- 62
"00001000000000000111001100001000", -- 63
"00000110110000100001000000010010", -- 64
"01001000100001000010000100001000", -- 65
"00000111000000000000000000000000", -- 66

-- ROM then filled with zero
    others => (others => '0'));
begin
  data <= Prom_ROM(conv_integer(unsigned(addr)));
end arch; 
